/*~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~*/ 
/*~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~*/
/* Engineer    : Lqc                                                         
/* File        : single_bit_s2f.v                                                         
/* Create      : 2022-08-29 20:54:12
/* Revise      : 2022-08-29 20:54:12                                                  
/* Module Name : single_bit_s2f                                                 
/* Description : 跨时钟域处理
/*               单比特信号慢时钟到快时钟处理方法
/*               边沿检测同步器      
/*  慢时钟域下的单比特信号的脉冲宽度，必须要大于或等于快时钟域下2个时钟
/*  周期。这样才能保证慢时钟域的脉冲信号是足够保持到被快时钟域的同步器拿到。                                                        
/* Editor : sublime text3, tab size (4)                                                                                
/*~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~*/
/*~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~*/

module single_bit_s2f(
	input         clka,         //slow clk
	input         clkb,         //fast clk
	input         rst,
	input         din,
	output        dout
	);

reg               din_reg1;
reg               din_reg2;
/*~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~*/
/*      Main Code                                                                  */
/*~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~*/
//在快时钟下对输入的信号打两拍做同步
always @(posedge clkb or posedge rst) begin
	if (rst) begin
		din_reg1 <= 'd0;
		din_reg2 <= 'd0;
	end
	else begin
		din_reg1 <= din;
		din_reg2 <= din_reg1;		
	end
end

//对打拍的信号生成在快时钟下的脉冲信号
assign dout = (din_reg1 & (~din_reg2));

endmodule